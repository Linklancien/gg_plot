module plot

import gg
import arrays { max, min }

// render_graph creat a graph at x, y with a width of w and an height of h
pub fn render_raw_graph(ctx gg.Context, x f32, y f32, w f32, h f32, abscice []f32, value []f32, name string) {
	max := max(value) or { panic('No max value') }
	min := min(value) or { panic('No min value') }
	max_a := max(abscice) or { panic('No max abscice') }

	f := fn [max, min, y, h] (value f32) f32 {
		return y + h - h * (value - min) / (max - min)
	}

	mut render_max := true
	mut render_min := true
	// Some magic numbers
	ctx.draw_rounded_rect_filled(f32(x - 10), f32(y - 10), f32(w + 35), f32(h + 10 + 35),
		5, gg.dark_gray)
	for k in 0 .. (abscice.len - 1) {
		ctx.draw_line(f32(x + w * abscice[k] / max_a), f32(f(value[k])), f32(x + w * abscice[k +
			1] / max_a), f32(f(value[k + 1])), gg.red)
		if k == 0 || k == abscice.len - 2 {
			ctx.draw_text_def(int(x + w * abscice[k] / max_a), int(f(value[k])), 'x: ${abscice[k]}  y: ${value[k]}')
			if value[k] == min {
				render_min = false
			}
			if value[k] == max {
				render_max = false
			}
		} else if value[k] == max && render_max {
			ctx.draw_text_def(int(x + w * abscice[k] / max_a), int(f(value[k])), 'x: ${abscice[k]}  y: ${value[k]}')
			render_max = false
		} else if value[k] == min && render_min {
			ctx.draw_text_def(int(x + w * abscice[k] / max_a), int(f(value[k])), 'x: ${abscice[k]}  y: ${value[k]}')
			render_min = false
		}
	}
	// ctx.draw_text_def(int(x), int(f(value[0])), '${value[0]}')
	// ctx.draw_text_def(int(x + w), int(f(value[abscice.len - 1])), '${value[abscice.len - 1]}')
	ctx.draw_text_def(int(x + w / 2), int(y + h + 10), name)
}

// utility
pub fn linear_interpolation(a f32, b f32, k f32, n f32) f32 {
	return a + (b - a) * k / n
}

//
// a: global position
// b: value the will be plot
// c: visuals
pub struct Diagram {
mut:
	// a:
	pos  Pos
	size Pos = Pos{x: 10, y: 10}

	// b:
	abscises [][]f32
	values   [][]f32
	colors   []gg.Color
	layers   []int

	// c:
	grid       Grid
	background gg.Color = gg.dark_gray
	border     f32      = 10
	corner     f32      = 5
	title      Label
	x_label    Label
	y_label    Label
}

struct Pos {
	x f32
	y f32
}

struct Label {
mut:
	text string
	cfg  gg.TextCfg
}

struct Grid {
	color gg.Color = gg.black
	x     bool     = true
	x_nb  int      = 5
	y     bool     = true
	y_nb  int      = 5
}

// creation
// basic creation
pub fn plot(abscises [][]f32, values [][]f32, colors []gg.Color, layers []int) Diagram {
	assert abscises.len == values.len, "Len of abscises and values doesn't match"
	assert abscises.len == colors.len, "Len of abscises and colors doesn't match"
	assert abscises.len == layers.len, "Len of abscises and layers doesn't match"
	return Diagram{
		abscises: abscises
		values:   values
		colors:   colors
		layers:	layers
	}
}

// changes
pub fn (mut dia Diagram) change_pos(x f32, y f32) {
	dia.pos = Pos{
		x: x
		y: y
	}
}

pub fn (mut dia Diagram) change_size(w f32, h f32) {
	dia.size = Pos{
		x: w
		y: h
	}
}

pub fn (mut dia Diagram) add_curve(abscice []f32, value []f32, color gg.Color, layer int) {
	dia.abscises << abscice
	dia.values << value
	dia.colors << color
	dia.layers << layer
}

pub fn (mut dia Diagram) show_grid(to_show bool) {
	dia.grid = Grid{
		x: to_show
		y: to_show
	}
}

pub fn (mut dia Diagram) title(text string) {
	dia.title.text = text
}

pub fn (mut dia Diagram) x_label(text string) {
	dia.x_label.text = text
}

pub fn (mut dia Diagram) y_label(text string) {
	dia.y_label.text = text
}

pub fn (mut dia Diagram) border_size(border f32) {
	dia.border = border
}

// rendering
pub fn (dia Diagram) render(ctx gg.Context) {
	// draw back
	ctx.draw_rounded_rect_filled(dia.pos.x, dia.pos.y, dia.size.x, dia.size.y, dia.corner,
		dia.background)
	// draw grid
	if dia.grid.x {
		dia.render_x_grid(ctx)
	}
	if dia.grid.y {
		dia.render_y_grid(ctx)
	}
	// draw curves
	max_x := dia.pos.x + dia.size.x - dia.border
	min_x := dia.pos.x + dia.border

	max_y := dia.pos.y + dia.size.y - dia.border
	min_y := dia.pos.y + dia.border

	list_max := dia.get_list_max()
	
	for id in 0 .. dia.abscises.len {
		render_curve(ctx, min_x, max_x, min_y, max_y, dia.abscises[id], dia.values[id],
			dia.colors[id], list_max[dia.layers[id]])
	}
	// draw axes

	// draw labels
}

// draw grid
fn (dia Diagram) render_x_grid(ctx gg.Context) {
	max_x := dia.pos.x + dia.size.x - dia.border
	min_x := dia.pos.x + dia.border

	max_y := dia.pos.y + dia.size.y - dia.border
	min_y := dia.pos.y + dia.border

	total := dia.grid.x_nb

	f := fn [min_x, max_x, total] (value f32) f32 {
		return linear_interpolation(min_x, max_x, value, total)
	}

	for i in 0 .. (total + 1) {
		x := f(i)
		ctx.draw_line(x, min_y, x, max_y, dia.grid.color)
	}
}

fn (dia Diagram) render_y_grid(ctx gg.Context) {
	max_x := dia.pos.x + dia.size.x - dia.border
	min_x := dia.pos.x + dia.border

	max_y := dia.pos.y + dia.size.y - dia.border
	min_y := dia.pos.y + dia.border

	total := dia.grid.x_nb

	f := fn [min_y, max_y, total] (value f32) f32 {
		return linear_interpolation(min_y, max_y, value, total)
	}

	for i in 0 .. (total + 1) {
		y := f(i)
		ctx.draw_line(min_x, y, max_x, y, dia.grid.color)
	}
}

// draw curves
fn (dia Diagram) get_list_max() []f32 {
	mut list_max := []f32{len: dia.values.len, init: max(dia.values[index]) or {panic('No max value for dia: $dia')}}
	for i, layer in dia.layers{
		max := max(dia.values[i]) or {panic('No max value for dia: $dia')}
		if list_max[layer] < max{
			list_max[layer] = max
		}
	}
	return list_max
}

fn render_curve(ctx gg.Context, min_x f32, max_x f32, min_y f32, max_y f32, abscice []f32, value []f32, color gg.Color, max_value f32) {
	max_abs := max(abscice) or { panic('no max abs') }
	f_x := fn [min_x, max_x, max_abs] (abs f32) f32 {
		return linear_interpolation(min_x, max_x, abs, max_abs)
	}

	f_y := fn [min_y, max_y, max_value] (value f32) f32 {
		return linear_interpolation(max_y, min_y, value, max_value)
	}

	for k in 0 .. (abscice.len - 1) {
		x1 := f_x(abscice[k])
		x2 := f_x(abscice[k + 1])
		y1 := f_y(value[k])
		y2 := f_y(value[k + 1])
		ctx.draw_line(x1, y1, x2, y2, color)
	}
}
